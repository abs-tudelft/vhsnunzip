library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package vhsnunzip_pkg is

  type byte_array is array (natural range <>) of std_logic_vector(7 downto 0);

end package vhsnunzip_pkg;
